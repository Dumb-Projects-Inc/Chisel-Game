module TopModule (
    input  wire clock,     // 100 MHz input clock
    input  wire reset,         // Reset button (active high)

    output wire [3:0] io_vga_red,     // VGA red signal
    output wire [3:0] io_vga_green,   // VGA green signal
    output wire [3:0] io_vga_blue,    // VGA blue signal
    output wire io_vga_hsync,         // VGA hsync
    output wire io_vga_vsync          // VGA vsync
);

    // Wires for PLL
    wire clk25MHz;
    wire pll_locked;

    // PLL instantiation (generated by Clocking Wizard)
    clk_wiz_0 pll_inst (
        .clk_in1(clock),
        .reset(reset),
        .clk_out1(clk25MHz),
        .locked(pll_locked)
    );

    // Chisel-generated VGA controller
    VGAController vga (
        .clock(clk25MHz),        // Base clock domain (still needed)
        .reset(~pll_locked),      // Hold reset until PLL locks
        .io_red(io_vga_red),
        .io_green(io_vga_green),
        .io_blue(io_vga_blue),
        .io_hsync(io_vga_hsync),
        .io_vsync(io_vga_vsync)
    );


endmodule